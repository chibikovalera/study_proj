module tb;

reg clk;
reg [255:0] pixel_vector;
wire [7:0] neuron_out;

// Подключаем main модуль
main uut (
    .clk(clk),
    .pixel_vector(pixel_vector),
    .neuron_out(neuron_out)
);

// Генератор тактового сигнала
initial begin
    clk = 0;
    forever #5 clk = ~clk; // период 10нс
end

// Задаем все 8 стрелок как маски
localparam [255:0] ARROW_UP = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000100000000,16'b0000001110000000,
    16'b0000011111000000,16'b0000111111100000,16'b0001111111110000,16'b0000000100000000,
    16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,
    16'b0000000100000000,16'b0000000100000000,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_UPLEFT = {
    16'b0000000000000000,16'b0000000000000000,16'b0011111110000000,16'b0011111100000000,
    16'b0011111000000000,16'b0011110000000000,16'b0011101000000000,16'b0011000100000000,
    16'b0010000010000000,16'b0000000001000000,16'b0000000000100000,16'b0000000000010000,
    16'b0000000000001000,16'b0000000000000100,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_LEFTDOWN = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000100,16'b0000000000001000,
    16'b0000000000010000,16'b0000000000100000,16'b0000000001000000,16'b0010000010000000,
    16'b0011000100000000,16'b0011101000000000,16'b0011110000000000,16'b0011111000000000,
    16'b0011111100000000,16'b0011111110000000,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_LEFT = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000001000000000,
    16'b0000011000000000,16'b0000111000000000,16'b0001111000000000,16'b0011111111111100,
    16'b0001111000000000,16'b0000111000000000,16'b0000011000000000,16'b0000001000000000,
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_DOWN = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000100000000,16'b0000000100000000,
    16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,
    16'b0000000100000000,16'b0001111111110000,16'b0000111111100000,16'b0000011111000000,
    16'b0000001110000000,16'b0000000100000000,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_UPRIGHT = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000111111100,16'b0000000011111100,
    16'b0000000001111100,16'b0000000000111100,16'b0000000001011100,16'b0000000010001100,
    16'b0000000100000100,16'b0000001000000000,16'b0000010000000000,16'b0000100000000000,
    16'b0001000000000000,16'b0010000000000000,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_DOWNRIGHT = {
    16'b0000000000000000,16'b0000000000000000,16'b0010000000000000,16'b0001000000000000,
    16'b0000100000000000,16'b0000010000000000,16'b0000001000000000,16'b0000000100000100,
    16'b0000000010001100,16'b0000000001011100,16'b0000000000111100,16'b0000000001111100,
    16'b0000000011111100,16'b0000000111111100,16'b0000000000000000,16'b0000000000000000
};

localparam [255:0] ARROW_RIGHT = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000000001000000,
    16'b0000000001100000,16'b0000000001110000,16'b0000000001111000,16'b0011111111111100,
    16'b0000000001111000,16'b0000000001110000,16'b0000000001100000,16'b0000000001000000,
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000000000000000
};

// Массив всех стрелок
reg [255:0] arrow_masks [0:7];
initial begin
    arrow_masks[0] = ARROW_UP;
    arrow_masks[1] = ARROW_UPLEFT;
    arrow_masks[2] = ARROW_LEFTDOWN;
    arrow_masks[3] = ARROW_LEFT;
    arrow_masks[4] = ARROW_DOWN;
    arrow_masks[5] = ARROW_UPRIGHT;
    arrow_masks[6] = ARROW_DOWNRIGHT;
    arrow_masks[7] = ARROW_RIGHT;
end

integer i;
reg [7:0] out_tmp;
initial begin
    for (i = 0; i < 8; i = i + 1) begin
        pixel_vector = arrow_masks[i];
        #30; // ждем обработку нейронами
        out_tmp = neuron_out;

        if (out_tmp == 8'b00000001)       $display("Arrow UP -> neuron_out = UP");
        else if (out_tmp == 8'b00000010)  $display("Arrow UPLEFT -> neuron_out = UPLEFT");
        else if (out_tmp == 8'b00000100)  $display("Arrow LEFTDOWN -> neuron_out = LEFTDOWN");
        else if (out_tmp == 8'b00001000)  $display("Arrow LEFT -> neuron_out = LEFT");
        else if (out_tmp == 8'b00010000)  $display("Arrow DOWN -> neuron_out = DOWN");
        else if (out_tmp == 8'b00100000)  $display("Arrow UPRIGHT -> neuron_out = UPRIGHT");
        else if (out_tmp == 8'b01000000)  $display("Arrow DOWNRIGHT -> neuron_out = DOWNRIGHT");
        else if (out_tmp == 8'b10000000)  $display("Arrow RIGHT -> neuron_out = RIGHT");
        else                               $display("Arrow UNKNOWN -> neuron_out = %b", out_tmp);

        #20;
    end

    $stop;
end

endmodule
