module main 
(
    input wire clk,
    input wire [255:0] pixel_vector,
    output wire [7:0] neuron_out
);

// 256-битные маски для нейронов
localparam [255:0] ARROW_UP = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000100000000,16'b0000001110000000,
    16'b0000011111000000,16'b0000111111100000,16'b0001111111110000,16'b0000000100000000,
    16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,
    16'b0000000100000000,16'b0000000100000000,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_UPLEFT = {
    16'b0000000000000000,16'b0000000000000000,16'b0011111110000000,16'b0011111100000000,
    16'b0011111000000000,16'b0011110000000000,16'b0011101000000000,16'b0011000100000000,
    16'b0010000010000000,16'b0000000001000000,16'b0000000000100000,16'b0000000000010000,
    16'b0000000000001000,16'b0000000000000100,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_LEFTDOWN = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000100,16'b0000000000001000,
    16'b0000000000010000,16'b0000000000100000,16'b0000000001000000,16'b0010000010000000,
    16'b0011000100000000,16'b0011101000000000,16'b0011110000000000,16'b0011111000000000,
    16'b0011111100000000,16'b0011111110000000,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_LEFT = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000001000000000,
    16'b0000011000000000,16'b0000111000000000,16'b0001111000000000,16'b0011111111111100,
    16'b0001111000000000,16'b0000111000000000,16'b0000011000000000,16'b0000001000000000,
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_DOWN = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000100000000,16'b0000000100000000,
    16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,16'b0000000100000000,
    16'b0000000100000000,16'b0001111111110000,16'b0000111111100000,16'b0000011111000000,
    16'b0000001110000000,16'b0000000100000000,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_UPRIGHT = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000111111100,16'b0000000011111100,
    16'b0000000001111100,16'b0000000000111100,16'b0000000001011100,16'b0000000010001100,
    16'b0000000100000100,16'b0000001000000000,16'b0000010000000000,16'b0000100000000000,
    16'b0001000000000000,16'b0010000000000000,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_DOWNRIGHT = {
    16'b0000000000000000,16'b0000000000000000,16'b0010000000000000,16'b0001000000000000,
    16'b0000100000000000,16'b0000010000000000,16'b0000001000000000,16'b0000000100000100,
    16'b0000000010001100,16'b0000000001011100,16'b0000000000111100,16'b0000000001111100,
    16'b0000000011111100,16'b0000000111111100,16'b0000000000000000,16'b0000000000000000
};
localparam [255:0] ARROW_RIGHT = {
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000000001000000,
    16'b0000000001100000,16'b0000000001110000,16'b0000000001111000,16'b0011111111111100,
    16'b0000000001111000,16'b0000000001110000,16'b0000000001100000,16'b0000000001000000,
    16'b0000000000000000,16'b0000000000000000,16'b0000000000000000,16'b0000000000000000
};

// Подключение нейронов
Neuron #(.k(ARROW_UP),        .b(32)) neuron0 (.x(pixel_vector), .clk(clk), .out(neuron_out[0]));
Neuron #(.k(ARROW_UPLEFT),    .b(36)) neuron1 (.x(pixel_vector), .clk(clk), .out(neuron_out[1]));
Neuron #(.k(ARROW_LEFTDOWN),  .b(36)) neuron2 (.x(pixel_vector), .clk(clk), .out(neuron_out[2]));
Neuron #(.k(ARROW_LEFT),      .b(32)) neuron3 (.x(pixel_vector), .clk(clk), .out(neuron_out[3]));
Neuron #(.k(ARROW_DOWN),      .b(32)) neuron4 (.x(pixel_vector), .clk(clk), .out(neuron_out[4]));
Neuron #(.k(ARROW_UPRIGHT),   .b(36)) neuron5 (.x(pixel_vector), .clk(clk), .out(neuron_out[5]));
Neuron #(.k(ARROW_DOWNRIGHT), .b(36)) neuron6 (.x(pixel_vector), .clk(clk), .out(neuron_out[6]));
Neuron #(.k(ARROW_RIGHT),     .b(32)) neuron7 (.x(pixel_vector), .clk(clk), .out(neuron_out[7]));

endmodule
